module add(a,b,out);
  input[16:0] a,b;
  output[16:0] out;
  assign out=a+b;
endmodule
